localparam
    Bgcolor = 12'h000,
    Fgcolor = 12'h3E7;
